`timescale 1ns/100ps

// -------------------------------- pre defined macros
import uvm_pkg::*;
`include "uvm_macros.svh"

// -------------------------------- UVM Environment YAPP Packet
`include "./yapp/yapp_packet.sv"

// --------------------------------------------------------- Sequences

// --------------------------------------------------------- Test cases
